module cglm

#include "@VROOT/external/cglm/src/affine.c"
#include "@VROOT/external/cglm/src/affine2d.c"
#include "@VROOT/external/cglm/src/bezier.c"
#include "@VROOT/external/cglm/src/box.c"
#include "@VROOT/external/cglm/src/cam.c"
#include "@VROOT/external/cglm/src/curve.c"
#include "@VROOT/external/cglm/src/ease.c"
#include "@VROOT/external/cglm/src/euler.c"
#include "@VROOT/external/cglm/src/frustum.c"
#include "@VROOT/external/cglm/src/io.c"
#include "@VROOT/external/cglm/src/ivec2.c"
#include "@VROOT/external/cglm/src/ivec3.c"
#include "@VROOT/external/cglm/src/ivec4.c"
#include "@VROOT/external/cglm/src/mat2.c"
#include "@VROOT/external/cglm/src/mat3.c"
#include "@VROOT/external/cglm/src/mat4.c"
#include "@VROOT/external/cglm/src/plane.c"
#include "@VROOT/external/cglm/src/project.c"
#include "@VROOT/external/cglm/src/quat.c"
#include "@VROOT/external/cglm/src/ray.c"
#include "@VROOT/external/cglm/src/sphere.c"
#include "@VROOT/external/cglm/src/vec2.c"
#include "@VROOT/external/cglm/src/vec3.c"
#include "@VROOT/external/cglm/src/vec4.c"
#include "@VROOT/external/cglm/src/clipspace/ortho_lh_no.c"
#include "@VROOT/external/cglm/src/clipspace/ortho_lh_zo.c"
#include "@VROOT/external/cglm/src/clipspace/ortho_rh_no.c"
#include "@VROOT/external/cglm/src/clipspace/ortho_rh_zo.c"
#include "@VROOT/external/cglm/src/clipspace/persp_lh_no.c"
#include "@VROOT/external/cglm/src/clipspace/persp_lh_zo.c"
#include "@VROOT/external/cglm/src/clipspace/persp_rh_no.c"
#include "@VROOT/external/cglm/src/clipspace/persp_rh_zo.c"
#include "@VROOT/external/cglm/src/clipspace/project_no.c"
#include "@VROOT/external/cglm/src/clipspace/project_zo.c"
#include "@VROOT/external/cglm/src/clipspace/view_lh_no.c"
#include "@VROOT/external/cglm/src/clipspace/view_lh_zo.c"
#include "@VROOT/external/cglm/src/clipspace/view_rh_no.c"
#include "@VROOT/external/cglm/src/clipspace/view_rh_zo.c"
