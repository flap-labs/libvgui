module main
import window

fn main() {
	win := window.create(1280, 720, "Testing VGUI")
	window.run()
	window.quit()
}
